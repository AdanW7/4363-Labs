parameter LW = 6'b100011 ; 
parameter SW = 6'b101011 ;
parameter no_op = 32'b0000000_0000000_0000000_0000000 ;
parameter ALUop = 6'b0 ;
parameter CINDC = 54 ;
parameter BEQINIT = 55 ;
//C:\Users\Kartik\Documents\solution_lab2_fall_2023\solution
string filename="/home/wodzi003/Downloads/handout/specific_tests/ALU/NAND/7/regs.dat";
string filename1="/home/wodzi003/Downloads/handout/specific_tests/ALU/NAND/7/dmem.dat";
string filename2="/home/wodzi003/Downloads/handout/specific_tests/ALU/NAND/7/imem.dat";
string filename3="/home/wodzi003/Downloads/handout/specific_tests/ALU/NAND/7/mem_result.dat";
string filename4="/home/wodzi003/Downloads/handout/specific_tests/ALU/NAND/7/regs_result.dat";
//string filename5="/home/wodzi003/Downloads/handout/specific_tests/ALU/NAND/7/pc_sequence.dat";